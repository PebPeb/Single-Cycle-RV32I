
//
//	datapath.v
//		RV32I datapath
//

// -------------------------------- //
//	By: Bryce Keen	
//	Created: 12/04/2022
// -------------------------------- //
//	Last Modified: 12/04/2022

// Change Log:	NA

module datapath();







endmodule





